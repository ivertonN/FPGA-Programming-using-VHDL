`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:29:44 05/24/2019 
// Design Name: 
// Module Name:    SumOneDigit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SumOneDigit(
    input [3:0] X_in,
    input [3:0] Y_in,
    input C_in,
    output C_out,
    output [3:0] Z_out
    );


endmodule
